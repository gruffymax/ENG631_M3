library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity T10_M3_clockDelayB is
    generic
    (
        g_cycles : integer  --
    );
    Port(
        i_sysClock : in STD_LOGIC;
        i_CE       : in STD_LOGIC
        );
end T10_M3_clockDelayB;

architecture archClockDelayB of T10_M3_clockDelayB is

begin
    
    
    
end archClockDelayB;