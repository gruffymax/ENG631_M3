--Team 10 - 762102 872403
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity T10_M3_segmentDecode is
    Port ( 
           i_BCDBuffer : in STD_LOGIC_VECTOR (3 downto 0);
           
           o_SegmentCathode : out STD_LOGIC_VECTOR (6 downto 0)
           );
end T10_M3_segmentDecode;

architecture archSegmentDecode of T10_M3_segmentDecode is
    
begin
with i_BCDBuffer select
    -- Cathodes are ACTIVE LOW
	o_SegmentCathode <=  "1000000" when "0000",  -- 0
	                     "1111001" when "0001",  -- 1
	                     "0100100" when "0010",  -- 2
	                     "0110000" when "0011",  -- 3
	                     "0011001" when "0100",  -- 4
	                     "0010010" when "0101",  -- 5
	                     "0000010" when "0110",  -- 6
	                     "1111000" when "0111",  -- 7
	                     "0000000" when "1000",  -- 8
	                     "0011000" when "1001",  -- 9
	                     "0001000" when "1010",  -- A
	                     "0000011" when "1011",  -- B
	                     "0100111" when "1100",  -- C
	                     "0100001" when "1101",  -- D
	                     "0000110" when "1110",  -- E
	                     "0001110" when "1111",  -- F
	                     "0000000" when others;

end archSegmentDecode;
